`timescale 1ns/1ns

module DataPath (clk,rst, regSrc, regDst, pcSrc, ALUSrc, ALUOp, regWrite, memWrite, memRead, flush, zero, opCode, func);
    input clk,rst;
endmodule